VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO 16b_FA
  CLASS BLOCK ;
  FOREIGN 16b_FA ;
  ORIGIN 0.000 0.000 ;
  SIZE 150.000 BY 340.000 ;
  PIN c15_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 90.420 11.870 93.150 12.145 ;
    END
  END c15_not
  PIN c15
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 83.070 9.795 93.150 10.130 ;
    END
  END c15
  PIN s5_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 134.480 229.350 137.210 229.625 ;
    END
  END s5_not
  PIN s5
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 127.130 227.275 137.210 227.610 ;
    END
  END s5
  PIN s0_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 134.500 327.985 137.230 328.260 ;
    END
  END s0_not
  PIN s0
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 127.150 325.910 137.230 326.245 ;
    END
  END s0
  PIN s6_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 134.480 209.380 137.210 209.655 ;
    END
  END s6_not
  PIN s6
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 127.130 207.305 137.210 207.640 ;
    END
  END s6
  PIN s1_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 134.300 308.260 137.030 308.535 ;
    END
  END s1_not
  PIN s1
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 126.950 306.185 137.030 306.520 ;
    END
  END s1
  PIN s7_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 134.480 189.715 137.210 189.990 ;
    END
  END s7_not
  PIN s7
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 127.130 187.640 137.210 187.975 ;
    END
  END s7
  PIN s2_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 134.455 288.615 137.185 288.890 ;
    END
  END s2_not
  PIN s2
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 127.105 286.540 137.185 286.875 ;
    END
  END s2
  PIN s8_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 134.520 169.875 137.250 170.150 ;
    END
  END s8_not
  PIN s8
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 127.170 167.800 137.250 168.135 ;
    END
  END s8
  PIN s3_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 134.455 268.820 137.185 269.095 ;
    END
  END s3_not
  PIN s3
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 127.105 266.745 137.185 267.080 ;
    END
  END s3
  PIN s9_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 134.320 150.150 137.050 150.425 ;
    END
  END s9_not
  PIN s9
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 126.970 148.075 137.050 148.410 ;
    END
  END s9
  PIN s4_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 134.375 249.065 137.105 249.340 ;
    END
  END s4_not
  PIN s4
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 127.025 246.990 137.105 247.325 ;
    END
  END s4
  PIN s10_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 134.475 130.505 137.205 130.780 ;
    END
  END s10_not
  PIN s10
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 127.125 128.430 137.205 128.765 ;
    END
  END s10
  PIN s11_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 134.475 110.710 137.205 110.985 ;
    END
  END s11_not
  PIN s11
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 127.125 108.635 137.205 108.970 ;
    END
  END s11
  PIN s12_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 134.395 90.955 137.125 91.230 ;
    END
  END s12_not
  PIN s12
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 127.045 88.880 137.125 89.215 ;
    END
  END s12
  PIN s13_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 134.500 71.240 137.230 71.515 ;
    END
  END s13_not
  PIN s13
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 127.150 69.165 137.230 69.500 ;
    END
  END s13
  PIN s14_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 134.500 51.270 137.230 51.545 ;
    END
  END s14_not
  PIN s14
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 127.150 49.195 137.230 49.530 ;
    END
  END s14
  PIN s15_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 134.500 31.605 137.230 31.880 ;
    END
  END s15_not
  PIN s15
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 127.150 29.530 137.230 29.865 ;
    END
  END s15
  PIN z
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 77.445 12.170 86.040 12.470 ;
    END
  END z
  PIN z_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT 77.415 11.635 83.395 11.905 ;
    END
  END z_not
  PIN c0_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 135.915 329.745 139.135 330.045 ;
    END
  END c0_b
  PIN c0_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 132.970 329.000 140.695 329.300 ;
    END
  END c0_not_b
  PIN a0_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 121.715 334.615 137.450 335.025 ;
    END
  END a0_b
  PIN a0_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 122.310 333.835 137.440 334.290 ;
    END
  END a0_not_b
  PIN a1_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 121.515 314.890 137.250 315.300 ;
    END
  END a1_b
  PIN a1_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 122.110 314.110 137.240 314.565 ;
    END
  END a1_not_b
  PIN a2_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 121.670 295.245 137.405 295.655 ;
    END
  END a2_b
  PIN a2_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 122.265 294.465 137.395 294.920 ;
    END
  END a2_not_b
  PIN a3_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 121.670 275.450 137.405 275.860 ;
    END
  END a3_b
  PIN a3_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 122.265 274.670 137.395 275.125 ;
    END
  END a3_not_b
  PIN a4_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 121.590 255.695 137.325 256.105 ;
    END
  END a4_b
  PIN a4_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 122.185 254.915 137.315 255.370 ;
    END
  END a4_not_b
  PIN a5_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 121.695 235.980 137.430 236.390 ;
    END
  END a5_b
  PIN a5_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 122.290 235.200 137.420 235.655 ;
    END
  END a5_not_b
  PIN a6_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 121.695 216.010 137.430 216.420 ;
    END
  END a6_b
  PIN a6_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 122.290 215.230 137.420 215.685 ;
    END
  END a6_not_b
  PIN a7_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 121.695 196.345 137.430 196.755 ;
    END
  END a7_b
  PIN a7_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 122.290 195.565 137.420 196.020 ;
    END
  END a7_not_b
  PIN VDD
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 0.485 195.620 0.495 195.630 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 1.885 196.940 1.895 196.950 ;
    END
  END VSS
  PIN a3_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 7.615 269.820 10.120 270.115 ;
    END
  END a3_not_f
  PIN b3
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 7.620 269.105 10.135 269.400 ;
    END
  END b3
  PIN b3_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 7.655 268.475 10.120 268.770 ;
    END
  END b3_not
  PIN a4_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 7.525 250.845 9.985 251.150 ;
    END
  END a4_f
  PIN a4_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 7.485 250.110 9.990 250.405 ;
    END
  END a4_not_f
  PIN b4
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 7.490 249.395 10.005 249.690 ;
    END
  END b4
  PIN b4_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 7.525 248.765 9.990 249.060 ;
    END
  END b4_not
  PIN a5_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 7.655 231.085 10.115 231.390 ;
    END
  END a5_f
  PIN a5_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 7.615 230.350 10.120 230.645 ;
    END
  END a5_not_f
  PIN b5
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 7.620 229.635 10.135 229.930 ;
    END
  END b5
  PIN b5_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 7.655 229.005 10.120 229.300 ;
    END
  END b5_not
  PIN a6_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 7.605 211.275 10.065 211.580 ;
    END
  END a6_f
  PIN a6_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 7.565 210.540 10.070 210.835 ;
    END
  END a6_not_f
  PIN b6
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 7.570 209.825 10.085 210.120 ;
    END
  END b6
  PIN b6_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 7.605 209.195 10.070 209.490 ;
    END
  END b6_not
  PIN a7_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 7.575 191.480 10.035 191.785 ;
    END
  END a7_f
  PIN a7_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 7.535 190.745 10.040 191.040 ;
    END
  END a7_not_f
  PIN b7
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 7.540 190.030 10.055 190.325 ;
    END
  END b7
  PIN b7_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 7.575 189.400 10.040 189.695 ;
    END
  END b7_not
  PIN a0_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 7.705 329.795 10.165 330.100 ;
    END
  END a0_f
  PIN a0_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 7.665 329.060 10.170 329.355 ;
    END
  END a0_not_f
  PIN b0
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 7.670 328.345 10.185 328.640 ;
    END
  END b0
  PIN b0_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 7.705 327.715 10.170 328.010 ;
    END
  END b0_not
  PIN a1_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 7.660 310.105 10.120 310.410 ;
    END
  END a1_f
  PIN a1_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 7.620 309.370 10.125 309.665 ;
    END
  END a1_not_f
  PIN b1
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 7.625 308.655 10.140 308.950 ;
    END
  END b1
  PIN b1_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 7.660 308.025 10.125 308.320 ;
    END
  END b1_not
  PIN a2_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 7.850 290.395 10.310 290.700 ;
    END
  END a2_f
  PIN a2_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 7.810 289.660 10.315 289.955 ;
    END
  END a2_not_f
  PIN b2
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 7.815 288.945 10.330 289.240 ;
    END
  END b2
  PIN b2_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 7.850 288.315 10.315 288.610 ;
    END
  END b2_not
  PIN a3_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 7.655 270.555 10.115 270.860 ;
    END
  END a3_f
  PIN c0_f
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 4.750 326.640 25.095 326.935 ;
    END
  END c0_f
  PIN c0_f_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 4.570 325.775 25.680 326.070 ;
    END
  END c0_f_not
  PIN b12_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 7.545 90.655 10.010 90.950 ;
    END
  END b12_not
  PIN a13_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 7.675 72.975 10.135 73.280 ;
    END
  END a13_f
  PIN a13_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 7.635 72.240 10.140 72.535 ;
    END
  END a13_not_f
  PIN b13
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 7.640 71.525 10.155 71.820 ;
    END
  END b13
  PIN b13_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 7.675 70.895 10.140 71.190 ;
    END
  END b13_not
  PIN a14_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 7.625 53.165 10.085 53.470 ;
    END
  END a14_f
  PIN a14_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 7.585 52.430 10.090 52.725 ;
    END
  END a14_not_f
  PIN b14
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 7.590 51.715 10.105 52.010 ;
    END
  END b14
  PIN b14_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 7.625 51.085 10.090 51.380 ;
    END
  END b14_not
  PIN a15_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 7.595 33.370 10.055 33.675 ;
    END
  END a15_f
  PIN a15_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 7.555 32.635 10.060 32.930 ;
    END
  END a15_not_f
  PIN b15
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 7.560 31.920 10.075 32.215 ;
    END
  END b15
  PIN b15_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 7.595 31.290 10.060 31.585 ;
    END
  END b15_not
  PIN a8_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 7.725 171.685 10.185 171.990 ;
    END
  END a8_f
  PIN a8_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 7.685 170.950 10.190 171.245 ;
    END
  END a8_not_f
  PIN b8
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 7.690 170.235 10.205 170.530 ;
    END
  END b8
  PIN b8_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 7.725 169.605 10.190 169.900 ;
    END
  END b8_not
  PIN a9_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 7.680 151.995 10.140 152.300 ;
    END
  END a9_f
  PIN a9_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 7.640 151.260 10.145 151.555 ;
    END
  END a9_not_f
  PIN b9
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 7.645 150.545 10.160 150.840 ;
    END
  END b9
  PIN b9_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 7.680 149.915 10.145 150.210 ;
    END
  END b9_not
  PIN a10_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 7.870 132.285 10.330 132.590 ;
    END
  END a10_f
  PIN a10_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 7.830 131.550 10.335 131.845 ;
    END
  END a10_not_f
  PIN b10
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 7.835 130.835 10.350 131.130 ;
    END
  END b10
  PIN b10_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 7.870 130.205 10.335 130.500 ;
    END
  END b10_not
  PIN a11_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 7.675 112.445 10.135 112.750 ;
    END
  END a11_f
  PIN a11_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 7.635 111.710 10.140 112.005 ;
    END
  END a11_not_f
  PIN b11
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 7.640 110.995 10.155 111.290 ;
    END
  END b11
  PIN b11_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal3 ;
        RECT 7.675 110.365 10.140 110.660 ;
    END
  END b11_not
  PIN a12_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 7.545 92.735 10.005 93.040 ;
    END
  END a12_f
  PIN a12_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 7.505 92.000 10.010 92.295 ;
    END
  END a12_not_f
  PIN b12
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal3 ;
        RECT 7.510 91.285 10.025 91.580 ;
    END
  END b12
  PIN a8_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 121.735 176.505 137.470 176.915 ;
    END
  END a8_b
  PIN a10_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 122.285 136.355 137.415 136.810 ;
    END
  END a10_not_b
  PIN a11_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 121.690 117.340 137.425 117.750 ;
    END
  END a11_b
  PIN a11_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 122.285 116.560 137.415 117.015 ;
    END
  END a11_not_b
  PIN a12_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 121.610 97.585 137.345 97.995 ;
    END
  END a12_b
  PIN a12_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 122.205 96.805 137.335 97.260 ;
    END
  END a12_not_b
  PIN a13_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 121.715 77.870 137.450 78.280 ;
    END
  END a13_b
  PIN a13_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 122.310 77.090 137.440 77.545 ;
    END
  END a13_not_b
  PIN a14_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 121.715 57.900 137.450 58.310 ;
    END
  END a14_b
  PIN a14_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 122.310 57.120 137.440 57.575 ;
    END
  END a14_not_b
  PIN a15_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 121.715 38.235 137.450 38.645 ;
    END
  END a15_b
  PIN a15_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 122.310 37.455 137.440 37.910 ;
    END
  END a15_not_b
  PIN a8_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 122.330 175.725 137.460 176.180 ;
    END
  END a8_not_b
  PIN a9_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 121.535 156.780 137.270 157.190 ;
    END
  END a9_b
  PIN a9_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 122.130 156.000 137.260 156.455 ;
    END
  END a9_not_b
  PIN a10_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal3 ;
        RECT 121.690 137.135 137.425 137.545 ;
    END
  END a10_b
  OBS
      LAYER Nwell ;
        RECT 7.985 4.245 137.250 336.340 ;
      LAYER Metal1 ;
        RECT 8.415 330.345 140.715 336.340 ;
        RECT 8.415 329.600 135.615 330.345 ;
        RECT 139.435 329.600 140.715 330.345 ;
        RECT 8.415 328.700 132.670 329.600 ;
        RECT 8.415 328.560 140.715 328.700 ;
        RECT 8.415 327.685 134.200 328.560 ;
        RECT 137.530 327.685 140.715 328.560 ;
        RECT 8.415 326.545 140.715 327.685 ;
        RECT 8.415 325.610 126.850 326.545 ;
        RECT 137.530 325.610 140.715 326.545 ;
        RECT 8.415 308.835 140.715 325.610 ;
        RECT 8.415 307.960 134.000 308.835 ;
        RECT 137.330 307.960 140.715 308.835 ;
        RECT 8.415 306.820 140.715 307.960 ;
        RECT 8.415 305.885 126.650 306.820 ;
        RECT 137.330 305.885 140.715 306.820 ;
        RECT 8.415 289.190 140.715 305.885 ;
        RECT 8.415 288.315 134.155 289.190 ;
        RECT 137.485 288.315 140.715 289.190 ;
        RECT 8.415 287.175 140.715 288.315 ;
        RECT 8.415 286.240 126.805 287.175 ;
        RECT 137.485 286.240 140.715 287.175 ;
        RECT 8.415 269.395 140.715 286.240 ;
        RECT 8.415 268.520 134.155 269.395 ;
        RECT 137.485 268.520 140.715 269.395 ;
        RECT 8.415 267.380 140.715 268.520 ;
        RECT 8.415 266.445 126.805 267.380 ;
        RECT 137.485 266.445 140.715 267.380 ;
        RECT 8.415 249.640 140.715 266.445 ;
        RECT 8.415 248.765 134.075 249.640 ;
        RECT 137.405 248.765 140.715 249.640 ;
        RECT 8.415 247.625 140.715 248.765 ;
        RECT 8.415 246.690 126.725 247.625 ;
        RECT 137.405 246.690 140.715 247.625 ;
        RECT 8.415 229.925 140.715 246.690 ;
        RECT 8.415 229.050 134.180 229.925 ;
        RECT 137.510 229.050 140.715 229.925 ;
        RECT 8.415 227.910 140.715 229.050 ;
        RECT 8.415 226.975 126.830 227.910 ;
        RECT 137.510 226.975 140.715 227.910 ;
        RECT 8.415 209.955 140.715 226.975 ;
        RECT 8.415 209.080 134.180 209.955 ;
        RECT 137.510 209.080 140.715 209.955 ;
        RECT 8.415 207.940 140.715 209.080 ;
        RECT 8.415 207.005 126.830 207.940 ;
        RECT 137.510 207.005 140.715 207.940 ;
        RECT 8.415 190.290 140.715 207.005 ;
        RECT 8.415 189.415 134.180 190.290 ;
        RECT 137.510 189.415 140.715 190.290 ;
        RECT 8.415 188.275 140.715 189.415 ;
        RECT 8.415 187.340 126.830 188.275 ;
        RECT 137.510 187.340 140.715 188.275 ;
        RECT 8.415 170.450 140.715 187.340 ;
        RECT 8.415 169.575 134.220 170.450 ;
        RECT 137.550 169.575 140.715 170.450 ;
        RECT 8.415 168.435 140.715 169.575 ;
        RECT 8.415 167.500 126.870 168.435 ;
        RECT 137.550 167.500 140.715 168.435 ;
        RECT 8.415 150.725 140.715 167.500 ;
        RECT 8.415 149.850 134.020 150.725 ;
        RECT 137.350 149.850 140.715 150.725 ;
        RECT 8.415 148.710 140.715 149.850 ;
        RECT 8.415 147.775 126.670 148.710 ;
        RECT 137.350 147.775 140.715 148.710 ;
        RECT 8.415 131.080 140.715 147.775 ;
        RECT 8.415 130.205 134.175 131.080 ;
        RECT 137.505 130.205 140.715 131.080 ;
        RECT 8.415 129.065 140.715 130.205 ;
        RECT 8.415 128.130 126.825 129.065 ;
        RECT 137.505 128.130 140.715 129.065 ;
        RECT 8.415 111.285 140.715 128.130 ;
        RECT 8.415 110.410 134.175 111.285 ;
        RECT 137.505 110.410 140.715 111.285 ;
        RECT 8.415 109.270 140.715 110.410 ;
        RECT 8.415 108.335 126.825 109.270 ;
        RECT 137.505 108.335 140.715 109.270 ;
        RECT 8.415 91.530 140.715 108.335 ;
        RECT 8.415 90.655 134.095 91.530 ;
        RECT 137.425 90.655 140.715 91.530 ;
        RECT 8.415 89.515 140.715 90.655 ;
        RECT 8.415 88.580 126.745 89.515 ;
        RECT 137.425 88.580 140.715 89.515 ;
        RECT 8.415 71.815 140.715 88.580 ;
        RECT 8.415 70.940 134.200 71.815 ;
        RECT 137.530 70.940 140.715 71.815 ;
        RECT 8.415 69.800 140.715 70.940 ;
        RECT 8.415 68.865 126.850 69.800 ;
        RECT 137.530 68.865 140.715 69.800 ;
        RECT 8.415 51.845 140.715 68.865 ;
        RECT 8.415 50.970 134.200 51.845 ;
        RECT 137.530 50.970 140.715 51.845 ;
        RECT 8.415 49.830 140.715 50.970 ;
        RECT 8.415 48.895 126.850 49.830 ;
        RECT 137.530 48.895 140.715 49.830 ;
        RECT 8.415 32.180 140.715 48.895 ;
        RECT 8.415 31.305 134.200 32.180 ;
        RECT 137.530 31.305 140.715 32.180 ;
        RECT 8.415 30.165 140.715 31.305 ;
        RECT 8.415 29.230 126.850 30.165 ;
        RECT 137.530 29.230 140.715 30.165 ;
        RECT 8.415 12.770 140.715 29.230 ;
        RECT 8.415 12.205 77.145 12.770 ;
        RECT 86.340 12.445 140.715 12.770 ;
        RECT 8.415 11.335 77.115 12.205 ;
        RECT 86.340 11.870 90.120 12.445 ;
        RECT 83.695 11.570 90.120 11.870 ;
        RECT 93.450 11.570 140.715 12.445 ;
        RECT 83.695 11.335 140.715 11.570 ;
        RECT 8.415 10.430 140.715 11.335 ;
        RECT 8.415 9.495 82.770 10.430 ;
        RECT 93.450 9.495 140.715 10.430 ;
        RECT 8.415 4.245 140.715 9.495 ;
      LAYER Metal2 ;
        RECT 4.655 4.195 140.605 336.340 ;
      LAYER Metal3 ;
        RECT 4.390 334.315 121.415 335.025 ;
        RECT 137.750 334.315 141.320 335.025 ;
        RECT 4.390 333.535 122.010 334.315 ;
        RECT 137.740 333.535 141.320 334.315 ;
        RECT 4.390 330.400 141.320 333.535 ;
        RECT 4.390 329.655 7.405 330.400 ;
        RECT 10.465 329.655 141.320 330.400 ;
        RECT 4.390 328.760 7.365 329.655 ;
        RECT 10.470 328.940 141.320 329.655 ;
        RECT 4.390 328.045 7.370 328.760 ;
        RECT 10.485 328.045 141.320 328.940 ;
        RECT 4.390 327.415 7.405 328.045 ;
        RECT 10.470 327.415 141.320 328.045 ;
        RECT 4.390 327.235 141.320 327.415 ;
        RECT 4.390 326.370 4.450 327.235 ;
        RECT 25.395 326.370 141.320 327.235 ;
        RECT 25.980 325.475 141.320 326.370 ;
        RECT 4.390 315.600 141.320 325.475 ;
        RECT 4.390 314.590 121.215 315.600 ;
        RECT 137.550 314.590 141.320 315.600 ;
        RECT 4.390 313.810 121.810 314.590 ;
        RECT 137.540 313.810 141.320 314.590 ;
        RECT 4.390 310.710 141.320 313.810 ;
        RECT 4.390 309.965 7.360 310.710 ;
        RECT 10.420 309.965 141.320 310.710 ;
        RECT 4.390 309.070 7.320 309.965 ;
        RECT 10.425 309.250 141.320 309.965 ;
        RECT 4.390 308.355 7.325 309.070 ;
        RECT 10.440 308.355 141.320 309.250 ;
        RECT 4.390 307.725 7.360 308.355 ;
        RECT 10.425 307.725 141.320 308.355 ;
        RECT 4.390 295.955 141.320 307.725 ;
        RECT 4.390 294.945 121.370 295.955 ;
        RECT 137.705 294.945 141.320 295.955 ;
        RECT 4.390 294.165 121.965 294.945 ;
        RECT 137.695 294.165 141.320 294.945 ;
        RECT 4.390 291.000 141.320 294.165 ;
        RECT 4.390 290.255 7.550 291.000 ;
        RECT 10.610 290.255 141.320 291.000 ;
        RECT 4.390 289.360 7.510 290.255 ;
        RECT 10.615 289.540 141.320 290.255 ;
        RECT 4.390 288.645 7.515 289.360 ;
        RECT 10.630 288.645 141.320 289.540 ;
        RECT 4.390 288.015 7.550 288.645 ;
        RECT 10.615 288.015 141.320 288.645 ;
        RECT 4.390 276.160 141.320 288.015 ;
        RECT 4.390 275.150 121.370 276.160 ;
        RECT 137.705 275.150 141.320 276.160 ;
        RECT 4.390 274.370 121.965 275.150 ;
        RECT 137.695 274.370 141.320 275.150 ;
        RECT 4.390 271.160 141.320 274.370 ;
        RECT 4.390 270.415 7.355 271.160 ;
        RECT 10.415 270.415 141.320 271.160 ;
        RECT 4.390 269.520 7.315 270.415 ;
        RECT 10.420 269.700 141.320 270.415 ;
        RECT 4.390 268.805 7.320 269.520 ;
        RECT 10.435 268.805 141.320 269.700 ;
        RECT 4.390 268.175 7.355 268.805 ;
        RECT 10.420 268.175 141.320 268.805 ;
        RECT 4.390 256.405 141.320 268.175 ;
        RECT 4.390 255.395 121.290 256.405 ;
        RECT 137.625 255.395 141.320 256.405 ;
        RECT 4.390 254.615 121.885 255.395 ;
        RECT 137.615 254.615 141.320 255.395 ;
        RECT 4.390 251.450 141.320 254.615 ;
        RECT 4.390 250.705 7.225 251.450 ;
        RECT 10.285 250.705 141.320 251.450 ;
        RECT 4.390 249.810 7.185 250.705 ;
        RECT 10.290 249.990 141.320 250.705 ;
        RECT 4.390 249.095 7.190 249.810 ;
        RECT 10.305 249.095 141.320 249.990 ;
        RECT 4.390 248.465 7.225 249.095 ;
        RECT 10.290 248.465 141.320 249.095 ;
        RECT 4.390 236.690 141.320 248.465 ;
        RECT 4.390 235.680 121.395 236.690 ;
        RECT 137.730 235.680 141.320 236.690 ;
        RECT 4.390 234.900 121.990 235.680 ;
        RECT 137.720 234.900 141.320 235.680 ;
        RECT 4.390 231.690 141.320 234.900 ;
        RECT 4.390 230.945 7.355 231.690 ;
        RECT 10.415 230.945 141.320 231.690 ;
        RECT 4.390 230.050 7.315 230.945 ;
        RECT 10.420 230.230 141.320 230.945 ;
        RECT 4.390 229.335 7.320 230.050 ;
        RECT 10.435 229.335 141.320 230.230 ;
        RECT 4.390 228.705 7.355 229.335 ;
        RECT 10.420 228.705 141.320 229.335 ;
        RECT 4.390 216.720 141.320 228.705 ;
        RECT 4.390 215.710 121.395 216.720 ;
        RECT 137.730 215.710 141.320 216.720 ;
        RECT 4.390 214.930 121.990 215.710 ;
        RECT 137.720 214.930 141.320 215.710 ;
        RECT 4.390 211.880 141.320 214.930 ;
        RECT 4.390 211.135 7.305 211.880 ;
        RECT 10.365 211.135 141.320 211.880 ;
        RECT 4.390 210.240 7.265 211.135 ;
        RECT 10.370 210.420 141.320 211.135 ;
        RECT 4.390 209.525 7.270 210.240 ;
        RECT 10.385 209.525 141.320 210.420 ;
        RECT 4.390 208.895 7.305 209.525 ;
        RECT 10.370 208.895 141.320 209.525 ;
        RECT 4.390 197.055 141.320 208.895 ;
        RECT 4.390 196.045 121.395 197.055 ;
        RECT 137.730 196.045 141.320 197.055 ;
        RECT 4.390 195.265 121.990 196.045 ;
        RECT 137.720 195.265 141.320 196.045 ;
        RECT 4.390 192.085 141.320 195.265 ;
        RECT 4.390 191.340 7.275 192.085 ;
        RECT 10.335 191.340 141.320 192.085 ;
        RECT 4.390 190.445 7.235 191.340 ;
        RECT 10.340 190.625 141.320 191.340 ;
        RECT 4.390 189.730 7.240 190.445 ;
        RECT 10.355 189.730 141.320 190.625 ;
        RECT 4.390 189.100 7.275 189.730 ;
        RECT 10.340 189.100 141.320 189.730 ;
        RECT 4.390 177.215 141.320 189.100 ;
        RECT 4.390 176.205 121.435 177.215 ;
        RECT 137.770 176.205 141.320 177.215 ;
        RECT 4.390 175.425 122.030 176.205 ;
        RECT 137.760 175.425 141.320 176.205 ;
        RECT 4.390 172.290 141.320 175.425 ;
        RECT 4.390 171.545 7.425 172.290 ;
        RECT 10.485 171.545 141.320 172.290 ;
        RECT 4.390 170.650 7.385 171.545 ;
        RECT 10.490 170.830 141.320 171.545 ;
        RECT 4.390 169.935 7.390 170.650 ;
        RECT 10.505 169.935 141.320 170.830 ;
        RECT 4.390 169.305 7.425 169.935 ;
        RECT 10.490 169.305 141.320 169.935 ;
        RECT 4.390 157.490 141.320 169.305 ;
        RECT 4.390 156.480 121.235 157.490 ;
        RECT 137.570 156.480 141.320 157.490 ;
        RECT 4.390 155.700 121.830 156.480 ;
        RECT 137.560 155.700 141.320 156.480 ;
        RECT 4.390 152.600 141.320 155.700 ;
        RECT 4.390 151.855 7.380 152.600 ;
        RECT 10.440 151.855 141.320 152.600 ;
        RECT 4.390 150.960 7.340 151.855 ;
        RECT 10.445 151.140 141.320 151.855 ;
        RECT 4.390 150.245 7.345 150.960 ;
        RECT 10.460 150.245 141.320 151.140 ;
        RECT 4.390 149.615 7.380 150.245 ;
        RECT 10.445 149.615 141.320 150.245 ;
        RECT 4.390 137.845 141.320 149.615 ;
        RECT 4.390 136.835 121.390 137.845 ;
        RECT 137.725 136.835 141.320 137.845 ;
        RECT 4.390 136.055 121.985 136.835 ;
        RECT 137.715 136.055 141.320 136.835 ;
        RECT 4.390 132.890 141.320 136.055 ;
        RECT 4.390 132.145 7.570 132.890 ;
        RECT 10.630 132.145 141.320 132.890 ;
        RECT 4.390 131.250 7.530 132.145 ;
        RECT 10.635 131.430 141.320 132.145 ;
        RECT 4.390 130.535 7.535 131.250 ;
        RECT 10.650 130.535 141.320 131.430 ;
        RECT 4.390 129.905 7.570 130.535 ;
        RECT 10.635 129.905 141.320 130.535 ;
        RECT 4.390 118.050 141.320 129.905 ;
        RECT 4.390 117.040 121.390 118.050 ;
        RECT 137.725 117.040 141.320 118.050 ;
        RECT 4.390 116.260 121.985 117.040 ;
        RECT 137.715 116.260 141.320 117.040 ;
        RECT 4.390 113.050 141.320 116.260 ;
        RECT 4.390 112.305 7.375 113.050 ;
        RECT 10.435 112.305 141.320 113.050 ;
        RECT 4.390 111.410 7.335 112.305 ;
        RECT 10.440 111.590 141.320 112.305 ;
        RECT 4.390 110.695 7.340 111.410 ;
        RECT 10.455 110.695 141.320 111.590 ;
        RECT 4.390 110.065 7.375 110.695 ;
        RECT 10.440 110.065 141.320 110.695 ;
        RECT 4.390 98.295 141.320 110.065 ;
        RECT 4.390 97.285 121.310 98.295 ;
        RECT 137.645 97.285 141.320 98.295 ;
        RECT 4.390 96.505 121.905 97.285 ;
        RECT 137.635 96.505 141.320 97.285 ;
        RECT 4.390 93.340 141.320 96.505 ;
        RECT 4.390 92.595 7.245 93.340 ;
        RECT 10.305 92.595 141.320 93.340 ;
        RECT 4.390 91.700 7.205 92.595 ;
        RECT 10.310 91.880 141.320 92.595 ;
        RECT 4.390 90.985 7.210 91.700 ;
        RECT 10.325 90.985 141.320 91.880 ;
        RECT 4.390 90.355 7.245 90.985 ;
        RECT 10.310 90.355 141.320 90.985 ;
        RECT 4.390 78.580 141.320 90.355 ;
        RECT 4.390 77.570 121.415 78.580 ;
        RECT 137.750 77.570 141.320 78.580 ;
        RECT 4.390 76.790 122.010 77.570 ;
        RECT 137.740 76.790 141.320 77.570 ;
        RECT 4.390 73.580 141.320 76.790 ;
        RECT 4.390 72.835 7.375 73.580 ;
        RECT 10.435 72.835 141.320 73.580 ;
        RECT 4.390 71.940 7.335 72.835 ;
        RECT 10.440 72.120 141.320 72.835 ;
        RECT 4.390 71.225 7.340 71.940 ;
        RECT 10.455 71.225 141.320 72.120 ;
        RECT 4.390 70.595 7.375 71.225 ;
        RECT 10.440 70.595 141.320 71.225 ;
        RECT 4.390 58.610 141.320 70.595 ;
        RECT 4.390 57.600 121.415 58.610 ;
        RECT 137.750 57.600 141.320 58.610 ;
        RECT 4.390 56.820 122.010 57.600 ;
        RECT 137.740 56.820 141.320 57.600 ;
        RECT 4.390 53.770 141.320 56.820 ;
        RECT 4.390 53.025 7.325 53.770 ;
        RECT 10.385 53.025 141.320 53.770 ;
        RECT 4.390 52.130 7.285 53.025 ;
        RECT 10.390 52.310 141.320 53.025 ;
        RECT 4.390 51.415 7.290 52.130 ;
        RECT 10.405 51.415 141.320 52.310 ;
        RECT 4.390 50.785 7.325 51.415 ;
        RECT 10.390 50.785 141.320 51.415 ;
        RECT 4.390 38.945 141.320 50.785 ;
        RECT 4.390 37.935 121.415 38.945 ;
        RECT 137.750 37.935 141.320 38.945 ;
        RECT 4.390 37.155 122.010 37.935 ;
        RECT 137.740 37.155 141.320 37.935 ;
        RECT 4.390 33.975 141.320 37.155 ;
        RECT 4.390 33.230 7.295 33.975 ;
        RECT 10.355 33.230 141.320 33.975 ;
        RECT 4.390 32.335 7.255 33.230 ;
        RECT 10.360 32.515 141.320 33.230 ;
        RECT 4.390 31.620 7.260 32.335 ;
        RECT 10.375 31.620 141.320 32.515 ;
        RECT 4.390 30.990 7.295 31.620 ;
        RECT 10.360 30.990 141.320 31.620 ;
        RECT 4.390 25.410 141.320 30.990 ;
  END
END 16b_FA
END LIBRARY

